module SPFP_ALU(
	input logic [31:0] n1,
	input logic [31:0] n2,
	input logic [1:0] s,
	output logic [31:0] z	
	);

endmodule